library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	5610	)	,
(	5599	)	,
(	5588	)	,
(	5577	)	,
(	5566	)	,
(	5555	)	,
(	5544	)	,
(	5533	)	,
(	5522	)	,
(	5511	)	,
(	5500	)	,
(	5489	)	,
(	5478	)	,
(	5468	)	,
(	5457	)	,
(	5446	)	,
(	5435	)	,
(	5425	)	,
(	5414	)	,
(	5403	)	,
(	5393	)	,
(	5382	)	,
(	5371	)	,
(	5361	)	,
(	5350	)	,
(	5340	)	,
(	5329	)	,
(	5319	)	,
(	5308	)	,
(	5298	)	,
(	5287	)	,
(	5277	)	,
(	5266	)	,
(	5256	)	,
(	5246	)	,
(	5235	)	,
(	5225	)	,
(	5215	)	,
(	5204	)	,
(	5194	)	,
(	5184	)	,
(	5174	)	,
(	5163	)	,
(	5153	)	,
(	5143	)	,
(	5133	)	,
(	5123	)	,
(	5113	)	,
(	5103	)	,
(	5093	)	,
(	5083	)	,
(	5073	)	,
(	5063	)	,
(	5053	)	,
(	5043	)	,
(	5033	)	,
(	5023	)	,
(	5013	)	,
(	5003	)	,
(	4993	)	,
(	4983	)	,
(	4973	)	,
(	4964	)	,
(	4954	)	,
(	4944	)	,
(	4934	)	,
(	4924	)	,
(	4915	)	,
(	4905	)	,
(	4895	)	,
(	4886	)	,
(	4876	)	,
(	4866	)	,
(	4857	)	,
(	4847	)	,
(	4838	)	,
(	4828	)	,
(	4819	)	,
(	4809	)	,
(	4800	)	,
(	4790	)	,
(	4781	)	,
(	4771	)	,
(	4762	)	,
(	4753	)	,
(	4743	)	,
(	4734	)	,
(	4724	)	,
(	4715	)	,
(	4706	)	,
(	4697	)	,
(	4687	)	,
(	4678	)	,
(	4669	)	,
(	4660	)	,
(	4650	)	,
(	4641	)	,
(	4632	)	,
(	4623	)	,
(	4614	)	,
(	4605	)	,
(	4596	)	,
(	4587	)	,
(	4578	)	,
(	4569	)	,
(	4560	)	,
(	4551	)	,
(	4542	)	,
(	4533	)	,
(	4524	)	,
(	4515	)	,
(	4506	)	,
(	4497	)	,
(	4488	)	,
(	4479	)	,
(	4471	)	,
(	4462	)	,
(	4453	)	,
(	4444	)	,
(	4435	)	,
(	4427	)	,
(	4418	)	,
(	4409	)	,
(	4401	)	,
(	4392	)	,
(	4383	)	,
(	4375	)	,
(	4366	)	,
(	4358	)	,
(	4349	)	,
(	4340	)	,
(	4332	)	,
(	4323	)	,
(	4315	)	,
(	4306	)	,
(	4298	)	,
(	4289	)	,
(	4281	)	,
(	4273	)	,
(	4264	)	,
(	4256	)	,
(	4247	)	,
(	4239	)	,
(	4231	)	,
(	4222	)	,
(	4214	)	,
(	4206	)	,
(	4198	)	,
(	4189	)	,
(	4181	)	,
(	4173	)	,
(	4165	)	,
(	4157	)	,
(	4148	)	,
(	4140	)	,
(	4132	)	,
(	4124	)	,
(	4116	)	,
(	4108	)	,
(	4100	)	,
(	4092	)	,
(	4084	)	,
(	4076	)	,
(	4068	)	,
(	4060	)	,
(	4052	)	,
(	4044	)	,
(	4036	)	,
(	4028	)	,
(	4020	)	,
(	4012	)	,
(	4004	)	,
(	3997	)	,
(	3989	)	,
(	3981	)	,
(	3973	)	,
(	3965	)	,
(	3958	)	,
(	3950	)	,
(	3942	)	,
(	3934	)	,
(	3927	)	,
(	3919	)	,
(	3911	)	,
(	3904	)	,
(	3896	)	,
(	3889	)	,
(	3881	)	,
(	3873	)	,
(	3866	)	,
(	3858	)	,
(	3851	)	,
(	3843	)	,
(	3836	)	,
(	3828	)	,
(	3821	)	,
(	3813	)	,
(	3806	)	,
(	3798	)	,
(	3791	)	,
(	3784	)	,
(	3776	)	,
(	3769	)	,
(	3762	)	,
(	3754	)	,
(	3747	)	,
(	3740	)	,
(	3732	)	,
(	3725	)	,
(	3718	)	,
(	3711	)	,
(	3703	)	,
(	3696	)	,
(	3689	)	,
(	3682	)	,
(	3675	)	,
(	3668	)	,
(	3660	)	,
(	3653	)	,
(	3646	)	,
(	3639	)	,
(	3632	)	,
(	3625	)	,
(	3618	)	,
(	3611	)	,
(	3604	)	,
(	3597	)	,
(	3590	)	,
(	3583	)	,
(	3576	)	,
(	3569	)	,
(	3562	)	,
(	3555	)	,
(	3548	)	,
(	3542	)	,
(	3535	)	,
(	3528	)	,
(	3521	)	,
(	3514	)	,
(	3508	)	,
(	3501	)	,
(	3494	)	,
(	3487	)	,
(	3480	)	,
(	3474	)	,
(	3467	)	,
(	3460	)	,
(	3454	)	,
(	3447	)	,
(	3440	)	,
(	3434	)	,
(	3427	)	,
(	3421	)	,
(	3414	)	,
(	3407	)	,
(	3401	)	,
(	3394	)	,
(	3388	)	,
(	3381	)	,
(	3375	)	,
(	3368	)	,
(	3362	)	,
(	3355	)	,
(	3349	)	,
(	3342	)	,
(	3336	)	,
(	3330	)	,
(	3323	)	,
(	3317	)	,
(	3310	)	,
(	3304	)	,
(	3298	)	,
(	3291	)	,
(	3285	)	,
(	3279	)	,
(	3273	)	,
(	3266	)	,
(	3260	)	,
(	3254	)	,
(	3248	)	,
(	3241	)	,
(	3235	)	,
(	3229	)	,
(	3223	)	,
(	3217	)	,
(	3211	)	,
(	3204	)	,
(	3198	)	,
(	3192	)	,
(	3186	)	,
(	3180	)	,
(	3174	)	,
(	3168	)	,
(	3162	)	,
(	3156	)	,
(	3150	)	,
(	3144	)	,
(	3138	)	,
(	3132	)	,
(	3126	)	,
(	3120	)	,
(	3114	)	,
(	3108	)	,
(	3102	)	,
(	3096	)	,
(	3091	)	,
(	3085	)	,
(	3079	)	,
(	3073	)	,
(	3067	)	,
(	3061	)	,
(	3056	)	,
(	3050	)	,
(	3044	)	,
(	3038	)	,
(	3033	)	,
(	3027	)	,
(	3021	)	,
(	3015	)	,
(	3010	)	,
(	3004	)	,
(	2998	)	,
(	2993	)	,
(	2987	)	,
(	2982	)	,
(	2976	)	,
(	2970	)	,
(	2965	)	,
(	2959	)	,
(	2954	)	,
(	2948	)	,
(	2943	)	,
(	2937	)	,
(	2932	)	,
(	2926	)	,
(	2921	)	,
(	2915	)	,
(	2910	)	,
(	2904	)	,
(	2899	)	,
(	2893	)	,
(	2888	)	,
(	2882	)	,
(	2877	)	,
(	2872	)	,
(	2866	)	,
(	2861	)	,
(	2856	)	,
(	2850	)	,
(	2845	)	,
(	2840	)	,
(	2834	)	,
(	2829	)	,
(	2824	)	,
(	2819	)	,
(	2813	)	,
(	2808	)	,
(	2803	)	,
(	2798	)	,
(	2793	)	,
(	2787	)	,
(	2782	)	,
(	2777	)	,
(	2772	)	,
(	2767	)	,
(	2762	)	,
(	2757	)	,
(	2752	)	,
(	2746	)	,
(	2741	)	,
(	2736	)	,
(	2731	)	,
(	2726	)	,
(	2721	)	,
(	2716	)	,
(	2711	)	,
(	2706	)	,
(	2701	)	,
(	2696	)	,
(	2691	)	,
(	2686	)	,
(	2681	)	,
(	2677	)	,
(	2672	)	,
(	2667	)	,
(	2662	)	,
(	2657	)	,
(	2652	)	,
(	2647	)	,
(	2642	)	,
(	2638	)	,
(	2633	)	,
(	2628	)	,
(	2623	)	,
(	2618	)	,
(	2614	)	,
(	2609	)	,
(	2604	)	,
(	2599	)	,
(	2595	)	,
(	2590	)	,
(	2585	)	,
(	2581	)	,
(	2576	)	,
(	2571	)	,
(	2567	)	,
(	2562	)	,
(	2557	)	,
(	2553	)	,
(	2548	)	,
(	2543	)	,
(	2539	)	,
(	2534	)	,
(	2530	)	,
(	2525	)	,
(	2521	)	,
(	2516	)	,
(	2512	)	,
(	2507	)	,
(	2502	)	,
(	2498	)	,
(	2494	)	,
(	2489	)	,
(	2485	)	,
(	2480	)	,
(	2476	)	,
(	2471	)	,
(	2467	)	,
(	2462	)	,
(	2458	)	,
(	2454	)	,
(	2449	)	,
(	2445	)	,
(	2441	)	,
(	2436	)	,
(	2432	)	,
(	2427	)	,
(	2423	)	,
(	2419	)	,
(	2415	)	,
(	2410	)	,
(	2406	)	,
(	2402	)	,
(	2397	)	,
(	2393	)	,
(	2389	)	,
(	2385	)	,
(	2381	)	,
(	2376	)	,
(	2372	)	,
(	2368	)	,
(	2364	)	,
(	2360	)	,
(	2356	)	,
(	2351	)	,
(	2347	)	,
(	2343	)	,
(	2339	)	,
(	2335	)	,
(	2331	)	,
(	2327	)	,
(	2323	)	,
(	2319	)	,
(	2315	)	,
(	2310	)	,
(	2306	)	,
(	2302	)	,
(	2298	)	,
(	2294	)	,
(	2290	)	,
(	2286	)	,
(	2282	)	,
(	2278	)	,
(	2275	)	,
(	2271	)	,
(	2267	)	,
(	2263	)	,
(	2259	)	,
(	2255	)	,
(	2251	)	,
(	2247	)	,
(	2243	)	,
(	2239	)	,
(	2236	)	,
(	2232	)	,
(	2228	)	,
(	2224	)	,
(	2220	)	,
(	2216	)	,
(	2213	)	,
(	2209	)	,
(	2205	)	,
(	2201	)	,
(	2197	)	,
(	2194	)	,
(	2190	)	,
(	2186	)	,
(	2182	)	,
(	2179	)	,
(	2175	)	,
(	2171	)	,
(	2168	)	,
(	2164	)	,
(	2160	)	,
(	2157	)	,
(	2153	)	,
(	2149	)	,
(	2146	)	,
(	2142	)	,
(	2138	)	,
(	2135	)	,
(	2131	)	,
(	2128	)	,
(	2124	)	,
(	2120	)	,
(	2117	)	,
(	2113	)	,
(	2110	)	,
(	2106	)	,
(	2103	)	,
(	2099	)	,
(	2096	)	,
(	2092	)	,
(	2089	)	,
(	2085	)	,
(	2082	)	,
(	2078	)	,
(	2075	)	,
(	2071	)	,
(	2068	)	,
(	2064	)	,
(	2061	)	,
(	2058	)	,
(	2054	)	,
(	2051	)	,
(	2047	)	,
(	2044	)	,
(	2041	)	,
(	2037	)	,
(	2034	)	,
(	2031	)	,
(	2027	)	,
(	2024	)	,
(	2020	)	,
(	2017	)	,
(	2014	)	,
(	2011	)	,
(	2007	)	,
(	2004	)	,
(	2001	)	,
(	1997	)	,
(	1994	)	,
(	1991	)	,
(	1988	)	,
(	1984	)	,
(	1981	)	,
(	1978	)	,
(	1975	)	,
(	1972	)	,
(	1968	)	,
(	1965	)	,
(	1962	)	,
(	1959	)	,
(	1956	)	,
(	1953	)	,
(	1949	)	,
(	1946	)	,
(	1943	)	,
(	1940	)	,
(	1937	)	,
(	1934	)	,
(	1931	)	,
(	1928	)	,
(	1924	)	,
(	1921	)	,
(	1918	)	,
(	1915	)	,
(	1912	)	,
(	1909	)	,
(	1906	)	,
(	1903	)	,
(	1900	)	,
(	1897	)	,
(	1894	)	,
(	1891	)	,
(	1888	)	,
(	1885	)	,
(	1882	)	,
(	1879	)	,
(	1876	)	,
(	1873	)	,
(	1870	)	,
(	1867	)	,
(	1864	)	,
(	1861	)	,
(	1859	)	,
(	1856	)	,
(	1853	)	,
(	1850	)	,
(	1847	)	,
(	1844	)	,
(	1841	)	,
(	1838	)	,
(	1835	)	,
(	1833	)	,
(	1830	)	,
(	1827	)	,
(	1824	)	,
(	1821	)	,
(	1819	)	,
(	1816	)	,
(	1813	)	,
(	1810	)	,
(	1807	)	,
(	1805	)	,
(	1802	)	,
(	1799	)	,
(	1796	)	,
(	1793	)	,
(	1791	)	,
(	1788	)	,
(	1785	)	,
(	1783	)	,
(	1780	)	,
(	1777	)	,
(	1774	)	,
(	1772	)	,
(	1769	)	,
(	1766	)	,
(	1764	)	,
(	1761	)	,
(	1758	)	,
(	1756	)	,
(	1753	)	,
(	1750	)	,
(	1748	)	,
(	1745	)	,
(	1743	)	,
(	1740	)	,
(	1737	)	,
(	1735	)	,
(	1732	)	,
(	1730	)	,
(	1727	)	,
(	1724	)	,
(	1722	)	,
(	1719	)	,
(	1717	)	,
(	1714	)	,
(	1712	)	,
(	1709	)	,
(	1707	)	,
(	1704	)	,
(	1702	)	,
(	1699	)	,
(	1697	)	,
(	1694	)	,
(	1692	)	,
(	1689	)	,
(	1687	)	,
(	1684	)	,
(	1682	)	,
(	1679	)	,
(	1677	)	,
(	1674	)	,
(	1672	)	,
(	1669	)	,
(	1667	)	,
(	1665	)	,
(	1662	)	,
(	1660	)	,
(	1657	)	,
(	1655	)	,
(	1653	)	,
(	1650	)	,
(	1648	)	,
(	1645	)	,
(	1643	)	,
(	1641	)	,
(	1638	)	,
(	1636	)	,
(	1634	)	,
(	1631	)	,
(	1629	)	,
(	1627	)	,
(	1624	)	,
(	1622	)	,
(	1620	)	,
(	1617	)	,
(	1615	)	,
(	1613	)	,
(	1611	)	,
(	1608	)	,
(	1606	)	,
(	1604	)	,
(	1602	)	,
(	1599	)	,
(	1597	)	,
(	1595	)	,
(	1593	)	,
(	1590	)	,
(	1588	)	,
(	1586	)	,
(	1584	)	,
(	1581	)	,
(	1579	)	,
(	1577	)	,
(	1575	)	,
(	1573	)	,
(	1571	)	,
(	1568	)	,
(	1566	)	,
(	1564	)	,
(	1562	)	,
(	1560	)	,
(	1558	)	,
(	1555	)	,
(	1553	)	,
(	1551	)	,
(	1549	)	,
(	1547	)	,
(	1545	)	,
(	1543	)	,
(	1541	)	,
(	1539	)	,
(	1536	)	,
(	1534	)	,
(	1532	)	,
(	1530	)	,
(	1528	)	,
(	1526	)	,
(	1524	)	,
(	1522	)	,
(	1520	)	,
(	1518	)	,
(	1516	)	,
(	1514	)	,
(	1512	)	,
(	1510	)	,
(	1508	)	,
(	1506	)	,
(	1504	)	,
(	1502	)	,
(	1500	)	,
(	1498	)	,
(	1496	)	,
(	1494	)	,
(	1492	)	,
(	1490	)	,
(	1488	)	,
(	1486	)	,
(	1484	)	,
(	1482	)	,
(	1480	)	,
(	1478	)	,
(	1476	)	,
(	1474	)	,
(	1472	)	,
(	1470	)	,
(	1469	)	,
(	1467	)	,
(	1465	)	,
(	1463	)	,
(	1461	)	,
(	1459	)	,
(	1457	)	,
(	1455	)	,
(	1453	)	,
(	1452	)	,
(	1450	)	,
(	1448	)	,
(	1446	)	,
(	1444	)	,
(	1442	)	,
(	1440	)	,
(	1439	)	,
(	1437	)	,
(	1435	)	,
(	1433	)	,
(	1431	)	,
(	1429	)	,
(	1428	)	,
(	1426	)	,
(	1424	)	,
(	1422	)	,
(	1420	)	,
(	1419	)	,
(	1417	)	,
(	1415	)	,
(	1413	)	,
(	1412	)	,
(	1410	)	,
(	1408	)	,
(	1406	)	,
(	1405	)	,
(	1403	)	,
(	1401	)	,
(	1399	)	,
(	1398	)	,
(	1396	)	,
(	1394	)	,
(	1392	)	,
(	1391	)	,
(	1389	)	,
(	1387	)	,
(	1386	)	,
(	1384	)	,
(	1382	)	,
(	1380	)	,
(	1379	)	,
(	1377	)	,
(	1375	)	,
(	1374	)	,
(	1372	)	,
(	1370	)	,
(	1369	)	,
(	1367	)	,
(	1365	)	,
(	1364	)	,
(	1362	)	,
(	1361	)	,
(	1359	)	,
(	1357	)	,
(	1356	)	,
(	1354	)	,
(	1352	)	,
(	1351	)	,
(	1349	)	,
(	1348	)	,
(	1346	)	,
(	1344	)	,
(	1343	)	,
(	1341	)	,
(	1340	)	,
(	1338	)	,
(	1336	)	,
(	1335	)	,
(	1333	)	,
(	1332	)	,
(	1330	)	,
(	1329	)	,
(	1327	)	,
(	1325	)	,
(	1324	)	,
(	1322	)	,
(	1321	)	,
(	1319	)	,
(	1318	)	,
(	1316	)	,
(	1315	)	,
(	1313	)	,
(	1312	)	,
(	1310	)	,
(	1309	)	,
(	1307	)	,
(	1306	)	,
(	1304	)	,
(	1303	)	,
(	1301	)	,
(	1300	)	,
(	1298	)	,
(	1297	)	,
(	1295	)	,
(	1294	)	,
(	1292	)	,
(	1291	)	,
(	1289	)	,
(	1288	)	,
(	1286	)	,
(	1285	)	,
(	1283	)	,
(	1282	)	,
(	1281	)	,
(	1279	)	,
(	1278	)	,
(	1276	)	,
(	1275	)	,
(	1273	)	,
(	1272	)	,
(	1271	)	,
(	1269	)	,
(	1268	)	,
(	1266	)	,
(	1265	)	,
(	1263	)	,
(	1262	)	,
(	1261	)	,
(	1259	)	,
(	1258	)	,
(	1257	)	,
(	1255	)	,
(	1254	)	,
(	1252	)	,
(	1251	)	,
(	1250	)	,
(	1248	)	,
(	1247	)	,
(	1246	)	,
(	1244	)	,
(	1243	)	,
(	1241	)	,
(	1240	)	,
(	1239	)	,
(	1237	)	,
(	1236	)	,
(	1235	)	,
(	1233	)	,
(	1232	)	,
(	1231	)	,
(	1229	)	,
(	1228	)	,
(	1227	)	,
(	1226	)	,
(	1224	)	,
(	1223	)	,
(	1222	)	,
(	1220	)	,
(	1219	)	,
(	1218	)	,
(	1216	)	,
(	1215	)	,
(	1214	)	,
(	1213	)	,
(	1211	)	,
(	1210	)	,
(	1209	)	,
(	1207	)	,
(	1206	)	,
(	1205	)	,
(	1204	)	,
(	1202	)	,
(	1201	)	,
(	1200	)	,
(	1199	)	,
(	1197	)	,
(	1196	)	,
(	1195	)	,
(	1194	)	,
(	1192	)	,
(	1191	)	,
(	1190	)	,
(	1189	)	,
(	1187	)	,
(	1186	)	,
(	1185	)	,
(	1184	)	,
(	1183	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1178	)	,
(	1176	)	,
(	1175	)	,
(	1174	)	,
(	1173	)	,
(	1172	)	,
(	1171	)	,
(	1169	)	,
(	1168	)	,
(	1167	)	,
(	1166	)	,
(	1165	)	,
(	1163	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1159	)	,
(	1158	)	,
(	1156	)	,
(	1155	)	,
(	1154	)	,
(	1153	)	,
(	1152	)	,
(	1151	)	,
(	1150	)	,
(	1148	)	,
(	1147	)	,
(	1146	)	,
(	1145	)	,
(	1144	)	,
(	1143	)	,
(	1142	)	,
(	1140	)	,
(	1139	)	,
(	1138	)	,
(	1137	)	,
(	1136	)	,
(	1135	)	,
(	1134	)	,
(	1133	)	,
(	1131	)	,
(	1130	)	,
(	1129	)	,
(	1128	)	,
(	1127	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1121	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1116	)	,
(	1115	)	,
(	1114	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1104	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1099	)	,
(	1098	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1090	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1080	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1068	)	,
(	1067	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1052	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1031	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1025	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1020	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	996	)	,
(	996	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	989	)	,
(	989	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	984	)	,
(	983	)	,
(	983	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	977	)	,
(	977	)	,
(	976	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	972	)	,
(	972	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	968	)	,
(	967	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	962	)	,
(	962	)	,
(	961	)	,
(	960	)	,
(	959	)	,
(	958	)	,
(	957	)	,
(	957	)	,
(	956	)	,
(	955	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	952	)	,
(	951	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	948	)	,
(	947	)	,
(	946	)	,
(	945	)	,
(	944	)	,
(	943	)	,
(	943	)	,
(	942	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	939	)	,
(	938	)	,
(	937	)	,
(	936	)	,
(	935	)	,
(	935	)	,
(	934	)	,
(	933	)	,
(	932	)	,
(	931	)	,
(	931	)	,
(	930	)	,
(	929	)	,
(	928	)	,
(	927	)	,
(	927	)	,
(	926	)	,
(	925	)	,
(	924	)	,
(	923	)	,
(	923	)	,
(	922	)	,
(	921	)	,
(	920	)	,
(	920	)	,
(	919	)	,
(	918	)	,
(	917	)	,
(	916	)	,
(	916	)	,
(	915	)	,
(	914	)	,
(	913	)	,
(	912	)	,
(	912	)	,
(	911	)	,
(	910	)	,
(	909	)	,
(	909	)	,
(	908	)	,
(	907	)	,
(	906	)	,
(	905	)	,
(	905	)	,
(	904	)	,
(	903	)	,
(	902	)	,
(	902	)	,
(	901	)	,
(	900	)	,
(	899	)	,
(	899	)	,
(	898	)	,
(	897	)	,
(	896	)	,
(	895	)	,
(	895	)	,
(	894	)	,
(	893	)	,
(	892	)	,
(	892	)	,
(	891	)	,
(	890	)	,
(	889	)	,
(	889	)	,
(	888	)	,
(	887	)	,
(	886	)	,
(	885	)	,
(	885	)	,
(	884	)	,
(	883	)	,
(	882	)	,
(	882	)	,
(	881	)	,
(	880	)	,
(	879	)	,
(	879	)	,
(	878	)	,
(	877	)	,
(	876	)	,
(	876	)	,
(	875	)	,
(	874	)	,
(	873	)	,
(	873	)	,
(	872	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	868	)	,
(	867	)	,
(	867	)	,
(	866	)	,
(	865	)	,
(	864	)	,
(	864	)	,
(	863	)	,
(	862	)	,
(	861	)	,
(	861	)	,
(	860	)	,
(	859	)	,
(	858	)	,
(	858	)	,
(	857	)	,
(	856	)	,
(	855	)	,
(	855	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	851	)	,
(	850	)	,
(	850	)	,
(	849	)	,
(	848	)	,
(	847	)	,
(	847	)	,
(	846	)	,
(	845	)	,
(	844	)	,
(	844	)	,
(	843	)	,
(	842	)	,
(	841	)	,
(	841	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	837	)	,
(	836	)	,
(	836	)	,
(	835	)	,
(	834	)	,
(	833	)	,
(	833	)	,
(	832	)	,
(	831	)	,
(	830	)	,
(	830	)	,
(	829	)	,
(	828	)	,
(	828	)	,
(	827	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	823	)	,
(	822	)	,
(	822	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	818	)	,
(	817	)	,
(	817	)	,
(	816	)	,
(	815	)	,
(	815	)	,
(	814	)	,
(	813	)	,
(	812	)	,
(	812	)	,
(	811	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	807	)	,
(	807	)	,
(	806	)	,
(	805	)	,
(	804	)	,
(	804	)	,
(	803	)	,
(	802	)	,
(	802	)	,
(	801	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	797	)	,
(	797	)	,
(	796	)	,
(	795	)	,
(	794	)	,
(	794	)	,
(	793	)	,
(	792	)	,
(	792	)	,
(	791	)	,
(	790	)	,
(	789	)	,
(	789	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	782	)	,
(	782	)	,
(	781	)	,
(	780	)	,
(	779	)	,
(	779	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	770	)	,
(	769	)	,
(	769	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	756	)	,
(	755	)	,
(	755	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	748	)	,
(	748	)	,
(	747	)	,
(	746	)	,
(	746	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	742	)	,
(	741	)	,
(	741	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	730	)	,
(	730	)	,
(	729	)	,
(	728	)	,
(	728	)	,
(	727	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	719	)	,
(	719	)	,
(	718	)	,
(	717	)	,
(	716	)	,
(	716	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	710	)	,
(	710	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	706	)	,
(	705	)	,
(	705	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	699	)	,
(	699	)	,
(	698	)	,
(	697	)	,
(	697	)	,
(	696	)	,
(	695	)	,
(	695	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	686	)	,
(	686	)	,
(	685	)	,
(	684	)	,
(	684	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	676	)	,
(	676	)	,
(	675	)	,
(	674	)	,
(	674	)	,
(	673	)	,
(	672	)	,
(	672	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	666	)	,
(	666	)	,
(	665	)	,
(	664	)	,
(	664	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	658	)	,
(	658	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	654	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	647	)	,
(	647	)	,
(	646	)	,
(	645	)	,
(	645	)	,
(	644	)	,
(	643	)	,
(	643	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	629	)	,
(	629	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	622	)	,
(	622	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	619	)	,
(	618	)	,
(	617	)	,
(	617	)	,
(	616	)	,
(	615	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	607	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	603	)	,
(	602	)	,
(	601	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	598	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	595	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	592	)	,
(	592	)	,
(	591	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	579	)	,
(	578	)	,
(	577	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	573	)	,
(	573	)	,
(	572	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	570	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	561	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	559	)	,
(	558	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	540	)	,
(	539	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	531	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	519	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	502	)	,
(	502	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	504	)	,
(	504	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	506	)	,
(	506	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	508	)	,
(	508	)	,
(	509	)	,
(	509	)	,
(	510	)	,
(	510	)	,
(	511	)	,
(	511	)	,
(	512	)	,
(	512	)	,
(	513	)	,
(	513	)	,
(	514	)	,
(	514	)	,
(	515	)	,
(	515	)	,
(	516	)	,
(	516	)	,
(	517	)	,
(	517	)	,
(	518	)	,
(	518	)	,
(	519	)	,
(	519	)	,
(	520	)	,
(	520	)	,
(	521	)	,
(	522	)	,
(	522	)	,
(	523	)	,
(	523	)	,
(	524	)	,
(	525	)	,
(	525	)	,
(	526	)	,
(	526	)	,
(	527	)	,
(	528	)	,
(	528	)	,
(	529	)	,
(	529	)	,
(	530	)	,
(	531	)	,
(	531	)	,
(	532	)	,
(	533	)	,
(	533	)	,
(	534	)	,
(	535	)	,
(	535	)	,
(	536	)	,
(	537	)	,
(	538	)	,
(	538	)	,
(	539	)	,
(	540	)	,
(	540	)	,
(	541	)	,
(	542	)	,
(	543	)	,
(	543	)	,
(	544	)	,
(	545	)	,
(	546	)	,
(	546	)	,
(	547	)	,
(	548	)	,
(	549	)	,
(	550	)	,
(	550	)	,
(	551	)	,
(	552	)	,
(	553	)	,
(	554	)	,
(	554	)	,
(	555	)	,
(	556	)	,
(	557	)	,
(	558	)	,
(	559	)	,
(	559	)	,
(	560	)	,
(	561	)	,
(	562	)	,
(	563	)	,
(	564	)	,
(	565	)	,
(	566	)	,
(	567	)	,
(	567	)	,
(	568	)	,
(	569	)	,
(	570	)	,
(	571	)	,
(	572	)	,
(	573	)	,
(	574	)	,
(	575	)	,
(	576	)	,
(	577	)	,
(	578	)	,
(	579	)	,
(	580	)	,
(	581	)	,
(	582	)	,
(	583	)	,
(	584	)	,
(	585	)	,
(	586	)	,
(	587	)	,
(	588	)	,
(	589	)	,
(	590	)	,
(	591	)	,
(	592	)	,
(	593	)	,
(	594	)	,
(	596	)	,
(	597	)	,
(	598	)	,
(	599	)	,
(	600	)	,
(	601	)	,
(	602	)	,
(	603	)	,
(	604	)	,
(	606	)	,
(	607	)	,
(	608	)	,
(	609	)	,
(	610	)	,
(	611	)	,
(	613	)	,
(	614	)	,
(	615	)	,
(	616	)	,
(	617	)	,
(	619	)	,
(	620	)	,
(	621	)	,
(	622	)	,
(	624	)	,
(	625	)	,
(	626	)	,
(	627	)	,
(	629	)	,
(	630	)	,
(	631	)	,
(	632	)	,
(	634	)	,
(	635	)	,
(	636	)	,
(	638	)	,
(	639	)	,
(	640	)	,
(	642	)	,
(	643	)	,
(	644	)	,
(	646	)	,
(	647	)	,
(	649	)	,
(	650	)	,
(	651	)	,
(	653	)	,
(	654	)	,
(	656	)	,
(	657	)	,
(	658	)	,
(	660	)	,
(	661	)	,
(	663	)	,
(	664	)	,
(	666	)	,
(	667	)	,
(	669	)	,
(	670	)	,
(	672	)	,
(	673	)	,
(	675	)	,
(	676	)	,
(	678	)	,
(	679	)	,
(	681	)	,
(	682	)	,
(	684	)	,
(	685	)	,
(	687	)	,
(	688	)	,
(	690	)	,
(	692	)	,
(	693	)	,
(	695	)	,
(	696	)	,
(	698	)	,
(	700	)	,
(	701	)	,
(	703	)	,
(	705	)	,
(	706	)	,
(	708	)	,
(	710	)	,
(	711	)	,
(	713	)	,
(	715	)	,
(	716	)	,
(	718	)	,
(	720	)	,
(	722	)	,
(	723	)	,
(	725	)	,
(	727	)	,
(	729	)	,
(	730	)	,
(	732	)	,
(	734	)	,
(	736	)	,
(	738	)	,
(	739	)	,
(	741	)	,
(	743	)	,
(	745	)	,
(	747	)	,
(	749	)	,
(	750	)	,
(	752	)	,
(	754	)	,
(	756	)	,
(	758	)	,
(	760	)	,
(	762	)	,
(	764	)	,
(	766	)	,
(	768	)	,
(	769	)	,
(	771	)	,
(	773	)	,
(	775	)	,
(	777	)	,
(	779	)	,
(	781	)	,
(	783	)	,
(	785	)	,
(	787	)	,
(	789	)	,
(	791	)	,
(	793	)	,
(	795	)	,
(	798	)	,
(	800	)	,
(	802	)	,
(	804	)	,
(	806	)	,
(	808	)	,
(	810	)	,
(	812	)	,
(	814	)	,
(	816	)	,
(	819	)	,
(	821	)	,
(	823	)	,
(	825	)	,
(	827	)	,
(	830	)	,
(	832	)	,
(	834	)	,
(	836	)	,
(	838	)	,
(	841	)	,
(	843	)	,
(	845	)	,
(	847	)	,
(	850	)	,
(	852	)	,
(	854	)	,
(	857	)	,
(	859	)	,
(	861	)	,
(	864	)	,
(	866	)	,
(	868	)	,
(	871	)	,
(	873	)	,
(	875	)	,
(	878	)	,
(	880	)	,
(	882	)	,
(	885	)	,
(	887	)	,
(	890	)	,
(	892	)	,
(	895	)	,
(	897	)	,
(	900	)	,
(	902	)	,
(	905	)	,
(	907	)	,
(	910	)	,
(	912	)	,
(	915	)	,
(	917	)	,
(	920	)	,
(	922	)	,
(	925	)	,
(	927	)	,
(	930	)	,
(	933	)	,
(	935	)	,
(	938	)	,
(	940	)	,
(	943	)	,
(	946	)	,
(	948	)	,
(	951	)	,
(	954	)	,
(	956	)	,
(	959	)	,
(	962	)	,
(	964	)	,
(	967	)	,
(	970	)	,
(	973	)	,
(	975	)	,
(	978	)	,
(	981	)	,
(	984	)	,
(	987	)	,
(	989	)	,
(	992	)	,
(	995	)	,
(	998	)	,
(	1001	)	,
(	1004	)	,
(	1006	)	,
(	1009	)	,
(	1012	)	,
(	1015	)	,
(	1018	)	,
(	1021	)	,
(	1024	)	,
(	1027	)	,
(	1030	)	,
(	1033	)	,
(	1036	)	,
(	1039	)	,
(	1042	)	,
(	1045	)	,
(	1048	)	,
(	1051	)	,
(	1054	)	,
(	1057	)	,
(	1060	)	,
(	1063	)	,
(	1066	)	,
(	1069	)	,
(	1072	)	,
(	1075	)	,
(	1078	)	,
(	1081	)	,
(	1085	)	,
(	1088	)	,
(	1091	)	,
(	1094	)	,
(	1097	)	,
(	1100	)	,
(	1104	)	,
(	1107	)	,
(	1110	)	,
(	1113	)	,
(	1117	)	,
(	1120	)	,
(	1123	)	,
(	1126	)	,
(	1130	)	,
(	1133	)	,
(	1136	)	,
(	1140	)	,
(	1143	)	,
(	1146	)	,
(	1150	)	,
(	1153	)	,
(	1156	)	,
(	1160	)	,
(	1163	)	,
(	1167	)	,
(	1170	)	,
(	1174	)	,
(	1177	)	,
(	1180	)	,
(	1184	)	,
(	1187	)	,
(	1191	)	,
(	1194	)	,
(	1198	)	,
(	1201	)	,
(	1205	)	,
(	1209	)	,
(	1212	)	,
(	1216	)	,
(	1219	)	,
(	1223	)	,
(	1227	)	,
(	1230	)	,
(	1234	)	,
(	1237	)	,
(	1241	)	,
(	1245	)	,
(	1248	)	,
(	1252	)	,
(	1256	)	,
(	1260	)	,
(	1263	)	,
(	1267	)	,
(	1271	)	,
(	1275	)	,
(	1278	)	,
(	1282	)	,
(	1286	)	,
(	1290	)	,
(	1294	)	,
(	1297	)	,
(	1301	)	,
(	1305	)	,
(	1309	)	,
(	1313	)	,
(	1317	)	,
(	1321	)	,
(	1325	)	,
(	1329	)	,
(	1333	)	,
(	1336	)	,
(	1340	)	,
(	1344	)	,
(	1348	)	,
(	1352	)	,
(	1356	)	,
(	1361	)	,
(	1365	)	,
(	1369	)	,
(	1373	)	,
(	1377	)	,
(	1381	)	,
(	1385	)	,
(	1389	)	,
(	1393	)	,
(	1397	)	,
(	1402	)	,
(	1406	)	,
(	1410	)	,
(	1414	)	,
(	1418	)	,
(	1423	)	,
(	1427	)	,
(	1431	)	,
(	1435	)	,
(	1440	)	,
(	1444	)	,
(	1448	)	,
(	1453	)	,
(	1457	)	,
(	1461	)	,
(	1466	)	,
(	1470	)	,
(	1474	)	,
(	1479	)	,
(	1483	)	,
(	1488	)	,
(	1492	)	,
(	1496	)	,
(	1501	)	,
(	1505	)	,
(	1510	)	,
(	1514	)	,
(	1519	)	,
(	1523	)	,
(	1528	)	,
(	1532	)	,
(	1537	)	,
(	1542	)	,
(	1546	)	,
(	1551	)	,
(	1555	)	,
(	1560	)	,
(	1565	)	,
(	1569	)	,
(	1574	)	,
(	1579	)	,
(	1583	)	,
(	1588	)	,
(	1593	)	,
(	1598	)	,
(	1602	)	,
(	1607	)	,
(	1612	)	,
(	1617	)	,
(	1622	)	,
(	1626	)	,
(	1631	)	,
(	1636	)	,
(	1641	)	,
(	1646	)	,
(	1651	)	,
(	1656	)	,
(	1661	)	,
(	1665	)	,
(	1670	)	,
(	1675	)	,
(	1680	)	,
(	1685	)	,
(	1690	)	,
(	1695	)	,
(	1700	)	,
(	1705	)	,
(	1711	)	,
(	1716	)	,
(	1721	)	,
(	1726	)	,
(	1731	)	,
(	1736	)	,
(	1741	)	,
(	1746	)	,
(	1752	)	,
(	1757	)	,
(	1762	)	,
(	1767	)	,
(	1772	)	,
(	1778	)	,
(	1783	)	,
(	1788	)	,
(	1794	)	,
(	1799	)	,
(	1804	)	,
(	1810	)	,
(	1815	)	,
(	1820	)	,
(	1826	)	,
(	1831	)	,
(	1836	)	,
(	1842	)	,
(	1847	)	,
(	1853	)	,
(	1858	)	,
(	1864	)	,
(	1869	)	,
(	1875	)	,
(	1880	)	,
(	1886	)	,
(	1891	)	,
(	1897	)	,
(	1903	)	,
(	1908	)	,
(	1914	)	,
(	1919	)	,
(	1925	)	,
(	1931	)	,
(	1936	)	,
(	1942	)	,
(	1948	)	,
(	1954	)	,
(	1959	)	,
(	1965	)	,
(	1971	)	,
(	1977	)	,
(	1982	)	,
(	1988	)	,
(	1994	)	,
(	2000	)	,
(	2006	)	,
(	2012	)	,
(	2018	)	,
(	2024	)	,
(	2030	)	,
(	2035	)	,
(	2041	)	,
(	2047	)	,
(	2053	)	,
(	2059	)	,
(	2065	)	,
(	2071	)	,
(	2078	)	,
(	2084	)	,
(	2090	)	,
(	2096	)	,
(	2102	)	,
(	2108	)	,
(	2114	)	,
(	2120	)	,
(	2127	)	,
(	2133	)	,
(	2139	)	,
(	2145	)	,
(	2151	)	,
(	2158	)	,
(	2164	)	,
(	2170	)	,
(	2177	)	,
(	2183	)	,
(	2189	)	,
(	2196	)	,
(	2202	)	,
(	2208	)	,
(	2215	)	,
(	2221	)	,
(	2228	)	,
(	2234	)	,
(	2241	)	,
(	2247	)	,
(	2254	)	,
(	2260	)	,
(	2267	)	,
(	2273	)	,
(	2280	)	,
(	2287	)	,
(	2293	)	,
(	2300	)	,
(	2306	)	,
(	2313	)	,
(	2320	)	,
(	2326	)	,
(	2333	)	,
(	2340	)	,
(	2347	)	,
(	2353	)	,
(	2360	)	,
(	2367	)	,
(	2374	)	,
(	2381	)	,
(	2387	)	,
(	2394	)	,
(	2401	)	,
(	2408	)	,
(	2415	)	,
(	2422	)	,
(	2429	)	,
(	2436	)	,
(	2443	)	,
(	2450	)	,
(	2457	)	,
(	2464	)	,
(	2471	)	,
(	2478	)	,
(	2485	)	,
(	2492	)	,
(	2499	)	,
(	2507	)	,
(	2514	)	,
(	2521	)	,
(	2528	)	,
(	2535	)	,
(	2543	)	,
(	2550	)	,
(	2557	)	,
(	2564	)	,
(	2572	)	,
(	2579	)	,
(	2586	)	,
(	2594	)	,
(	2601	)	,
(	2608	)	,
(	2616	)	,
(	2623	)	,
(	2631	)	,
(	2638	)	,
(	2646	)	,
(	2653	)	,
(	2661	)	,
(	2668	)	,
(	2676	)	,
(	2683	)	,
(	2691	)	,
(	2699	)	,
(	2706	)	,
(	2714	)	,
(	2722	)	,
(	2729	)	,
(	2737	)	,
(	2745	)	,
(	2752	)	,
(	2760	)	,
(	2768	)	,
(	2776	)	,
(	2783	)	,
(	2791	)	,
(	2799	)	,
(	2807	)	,
(	2815	)	,
(	2823	)	,
(	2831	)	,
(	2839	)	,
(	2847	)	,
(	2855	)	,
(	2863	)	,
(	2871	)	,
(	2879	)	,
(	2887	)	,
(	2895	)	,
(	2903	)	,
(	2911	)	,
(	2919	)	,
(	2927	)	,
(	2935	)	,
(	2944	)	,
(	2952	)	,
(	2960	)	,
(	2968	)	,
(	2977	)	,
(	2985	)	,
(	2993	)	,
(	3002	)	,
(	3010	)	,
(	3018	)	,
(	3027	)	,
(	3035	)	,
(	3043	)	,
(	3052	)	,
(	3060	)	,
(	3069	)	,
(	3077	)	,
(	3086	)	,
(	3094	)	,
(	3103	)	,
(	3111	)	,
(	3120	)	,
(	3129	)	,
(	3137	)	,
(	3146	)	,
(	3155	)	,
(	3163	)	,
(	3172	)	,
(	3181	)	,
(	3190	)	,
(	3198	)	,
(	3207	)	,
(	3216	)	,
(	3225	)	,
(	3234	)	,
(	3242	)	,
(	3251	)	,
(	3260	)	,
(	3269	)	,
(	3278	)	,
(	3287	)	,
(	3296	)	,
(	3305	)	,
(	3314	)	,
(	3323	)	,
(	3332	)	,
(	3341	)	,
(	3351	)	,
(	3360	)	,
(	3369	)	,
(	3378	)	,
(	3387	)	,
(	3396	)	,
(	3406	)	,
(	3415	)	,
(	3424	)	,
(	3434	)	,
(	3443	)	,
(	3452	)	,
(	3462	)	,
(	3471	)	,
(	3480	)	,
(	3490	)	,
(	3499	)	,
(	3509	)	,
(	3518	)	,
(	3528	)	,
(	3537	)	,
(	3547	)	,
(	3556	)	,
(	3566	)	,
(	3576	)	,
(	3585	)	,
(	3595	)	,
(	3605	)	,
(	3614	)	,
(	3624	)	,
(	3634	)	,
(	3643	)	,
(	3653	)	,
(	3663	)	,
(	3673	)	,
(	3683	)	,
(	3693	)	,
(	3702	)	,
(	3712	)	,
(	3722	)	,
(	3732	)	,
(	3742	)	,
(	3752	)	,
(	3762	)	,
(	3772	)	,
(	3782	)	,
(	3792	)	,
(	3803	)	,
(	3813	)	,
(	3823	)	,
(	3833	)	,
(	3843	)	,
(	3853	)	,
(	3864	)	,
(	3874	)	,
(	3884	)	,
(	3895	)	,
(	3905	)	,
(	3915	)	,
(	3926	)	,
(	3936	)	,
(	3946	)	,
(	3957	)	,
(	3967	)	,
(	3978	)	,
(	3988	)	,
(	3999	)	,
(	4009	)	,
(	4020	)	,
(	4031	)	,
(	4041	)	,
(	4052	)	,
(	4062	)	,
(	4073	)	,
(	4084	)	,
(	4095	)	,
(	4105	)	,
(	4116	)	,
(	4127	)	,
(	4138	)	,
(	4149	)	,
(	4159	)	,
(	4170	)	,
(	4181	)	,
(	4192	)	,
(	4203	)	,
(	4214	)	,
(	4225	)	,
(	4236	)	,
(	4247	)	,
(	4258	)	,
(	4269	)	,
(	4280	)	,
(	4292	)	,
(	4303	)	,
(	4314	)	,
(	4325	)	,
(	4336	)	,
(	4348	)	,
(	4359	)	,
(	4370	)	,
(	4382	)	,
(	4393	)	,
(	4404	)	,
(	4416	)	,
(	4427	)	,
(	4439	)	,
(	4450	)	,
(	4462	)	,
(	4473	)	,
(	4485	)	,
(	4496	)	,
(	4508	)	,
(	4519	)	,
(	4531	)	,
(	4543	)	,
(	4554	)	,
(	4566	)	,
(	4578	)	,
(	4590	)	,
(	4601	)	,
(	4613	)	,
(	4625	)	,
(	4637	)	,
(	4649	)	,
(	4661	)	,
(	4672	)	,
(	4684	)	,
(	4696	)	,
(	4708	)	,
(	4720	)	,
(	4732	)	,
(	4745	)	,
(	4757	)	,
(	4769	)	,
(	4781	)	,
(	4793	)	,
(	4805	)	,
(	4817	)	,
(	4830	)	,
(	4842	)	,
(	4854	)	,
(	4867	)	,
(	4879	)	,
(	4891	)	,
(	4904	)	,
(	4916	)	,
(	4929	)	,
(	4941	)	,
(	4953	)	,
(	4966	)	,
(	4979	)	,
(	4991	)	,
(	5004	)	,
(	5016	)	,
(	5029	)	,
(	5042	)	,
(	5054	)	,
(	5067	)	,
(	5080	)	,
(	5092	)	,
(	5105	)	,
(	5118	)	,
(	5131	)	,
(	5144	)	,
(	5157	)	,
(	5170	)	,
(	5183	)	,
(	5196	)	,
(	5208	)	,
(	5222	)	,
(	5235	)	,
(	5248	)	,
(	5261	)	,
(	5274	)	,
(	5287	)	,
(	5300	)	,
(	5313	)	,
(	5327	)	,
(	5340	)	,
(	5353	)	,
(	5366	)	,
(	5380	)	,
(	5393	)	,
(	5406	)	,
(	5420	)	,
(	5433	)	,
(	5447	)	,
(	5460	)	,
(	5474	)	,
(	5487	)	,
(	5501	)	,
(	5514	)	,
(	5528	)	,
(	5542	)	,
(	5555	)	,
(	5569	)	,
(	5583	)	,
(	5597	)	,
(	5610	)	,
(	5624	)	,
(	5638	)	,
(	5652	)	,
(	5666	)	,
(	5680	)	,
(	5693	)	,
(	5707	)	,
(	5721	)	,
(	5735	)	,
(	5749	)	,
(	5764	)	,
(	5778	)	,
(	5792	)	,
(	5806	)	,
(	5820	)	,
(	5834	)	,
(	5849	)	,
(	5863	)	,
(	5877	)	,
(	5891	)	,
(	5906	)	,
(	5920	)	,
(	5934	)	,
(	5949	)	,
(	5963	)	,
(	5978	)	,
(	5992	)	,
(	6007	)	,
(	6021	)	,
(	6036	)	,
(	6051	)	,
(	6065	)	,
(	6080	)	,
(	6095	)	,
(	6109	)	,
(	6124	)	,
(	6139	)	,
(	6154	)	,
(	6168	)	,
(	6183	)	,
(	6198	)	,
(	6213	)	,
(	6228	)	,
(	6243	)	,
(	6258	)	,
(	6273	)	,
(	6288	)	,
(	6303	)	,
(	6318	)	,
(	6333	)	,
(	6349	)	,
(	6364	)	,
(	6379	)	,
(	6394	)	,
(	6410	)	,
(	6425	)	,
(	6440	)	,
(	6456	)	,
(	6471	)	,
(	6486	)	,
(	6502	)	,
(	6517	)	,
(	6533	)	,
(	6548	)	,
(	6564	)	,
(	6580	)	,
(	6595	)	,
(	6611	)	,
(	6626	)	,
(	6642	)	,
(	6658	)	,
(	6674	)	,
(	6689	)	,
(	6705	)	,
(	6721	)	,
(	6737	)	,
(	6753	)	,
(	6769	)	,
(	6785	)	,
(	6801	)	,
(	6817	)	,
(	6833	)	,
(	6849	)	,
(	6865	)	,
(	6881	)	,
(	6897	)	,
(	6914	)	,
(	6930	)	,
(	6946	)	,
(	6962	)	,
(	6979	)	,
(	6995	)	,
(	7012	)	,
(	7028	)	,
(	7044	)	,
(	7061	)	,
(	7077	)	,
(	7094	)	,
(	7110	)	,
(	7127	)	,
(	7144	)	,
(	7160	)	,
(	7177	)	,
(	7194	)	,
(	7210	)	,
(	7227	)	,
(	7244	)	,
(	7261	)	,
(	7278	)	,
(	7295	)	,
(	7312	)	,
(	7328	)	,
(	7345	)	,
(	7362	)	,
(	7380	)	,
(	7397	)	,
(	7414	)	,
(	7431	)	,
(	7448	)	,
(	7465	)	,
(	7482	)	,
(	7500	)	,
(	7517	)	,
(	7534	)	,
(	7552	)	,
(	7569	)	,
(	7586	)	,
(	7604	)	,
(	7621	)	,
(	7639	)	,
(	7656	)	,
(	7674	)	,
(	7692	)	,
(	7709	)	,
(	7727	)	,
(	7744	)	,
(	7762	)	,
(	7780	)	,
(	7798	)	,
(	7816	)	,
(	7833	)	,
(	7851	)	,
(	7869	)	,
(	7887	)	,
(	7905	)	,
(	7923	)	,
(	7941	)	,
(	7959	)	,
(	7977	)	,
(	7995	)	,
(	8014	)	,
(	8032	)	,
(	8050	)	,
(	8068	)	,
(	8087	)	,
(	8105	)	,
(	8123	)	,
(	8142	)	,
(	8160	)	,
(	8178	)	,
(	8197	)	,
(	8215	)	,
(	8234	)	,
(	8253	)	,
(	8271	)	,
(	8290	)	,
(	8308	)	,
(	8327	)	,
(	8346	)	,
(	8365	)	,
(	8383	)	,
(	8402	)	,
(	8421	)	,
(	8440	)	,
(	8459	)	,
(	8478	)	,
(	8497	)	,
(	8516	)	,
(	8535	)	,
(	8554	)	,
(	8573	)	,
(	8592	)	,
(	8612	)	,
(	8631	)	,
(	8650	)	,
(	8669	)	,
(	8689	)	,
(	8708	)	,
(	8727	)	,
(	8747	)	,
(	8766	)	,
(	8786	)	,
(	8805	)	,
(	8825	)	,
(	8844	)	,
(	8864	)	,
(	8884	)	,
(	8903	)	,
(	8923	)	,
(	8943	)	,
(	8963	)	,
(	8983	)	,
(	9002	)	,
(	9022	)	,
(	9042	)	,
(	9062	)	,
(	9082	)	,
(	9102	)	,
(	9122	)	,
(	9142	)	,
(	9162	)	,
(	9183	)	,
(	9203	)	,
(	9223	)	,
(	9243	)	,
(	9264	)	,
(	9284	)	,
(	9304	)	,
(	9325	)	,
(	9345	)	,
(	9366	)	,
(	9386	)	,
(	9407	)	,
(	9427	)	,
(	9448	)	,
(	9468	)	,
(	9489	)	,
(	9510	)	,
(	9531	)	,
(	9551	)	,
(	9572	)	,
(	9593	)	,
(	9614	)	,
(	9635	)	,
(	9656	)	,
(	9677	)	,
(	9698	)	,
(	9719	)	,
(	9740	)	,
(	9761	)	,
(	9782	)	,
(	9803	)	,
(	9825	)	,
(	9846	)	,
(	9867	)	,
(	9888	)	,
(	9910	)	,
(	9931	)	,
(	9953	)	,
(	9974	)	,
(	9996	)	,
(	10017	)	,
(	10039	)	,
(	10060	)	,
(	10082	)	,
(	10104	)	,
(	10125	)	,
(	10147	)	,
(	10169	)	,
(	10191	)	,
(	10213	)	,
(	10235	)	,
(	10256	)	,
(	10278	)	,
(	10300	)	,
(	10322	)	,
(	10345	)	,
(	10367	)	,
(	10389	)	,
(	10411	)	,
(	10433	)	,
(	10456	)	,
(	10478	)	,
(	10500	)	,
(	10523	)	,
(	10545	)	,
(	10567	)	,
(	10590	)	,
(	10612	)	,
(	10635	)	,
(	10657	)	,
(	10680	)	,
(	10703	)	,
(	10725	)	,
(	10748	)	,
(	10771	)	,
(	10794	)	,
(	10817	)	,
(	10839	)	,
(	10862	)	,
(	10885	)	,
(	10908	)	,
(	10931	)	,
(	10954	)	,
(	10978	)	,
(	11001	)	,
(	11024	)	,
(	11047	)	,
(	11070	)	,
(	11094	)	,
(	11117	)	,
(	11140	)	,
(	11164	)	,
(	11187	)	,
(	11211	)	,
(	11234	)	,
(	11258	)	,
(	11281	)	,
(	11305	)	,
(	11329	)	,
(	11352	)	,
(	11376	)	,
(	11400	)	,
(	11424	)	,
(	11447	)	,
(	11471	)	,
(	11495	)	,
(	11519	)	,
(	11543	)	,
(	11567	)	,
(	11591	)	,
(	11615	)	,
(	11640	)	,
(	11664	)	,
(	11688	)	,
(	11712	)	,
(	11737	)	,
(	11761	)	,
(	11785	)	,
(	11810	)	,
(	11834	)	,
(	11859	)	,
(	11883	)	,
(	11908	)	,
(	11932	)	,
(	11957	)	,
(	11982	)	,
(	12006	)	,
(	12031	)	,
(	12056	)	,
(	12081	)	,
(	12106	)	,
(	12131	)	,
(	12156	)	,
(	12181	)	,
(	12206	)	,
(	12231	)	,
(	12256	)	,
(	12281	)	,
(	12306	)	,
(	12331	)	,
(	12357	)	,
(	12382	)	,
(	12407	)	,
(	12433	)	,
(	12458	)	,
(	12484	)	,
(	12509	)	,
(	12535	)	,
(	12560	)	,
(	12586	)	,
(	12612	)	,
(	12637	)	,
(	12663	)	,
(	12689	)	,
(	12715	)	,
(	12741	)	,
(	12766	)	,
(	12792	)	,
(	12818	)	,
(	12844	)	,
(	12870	)	,
(	12897	)	,
(	12923	)	,
(	12949	)	,
(	12975	)	,
(	13001	)	,
(	13028	)	,
(	13054	)	,
(	13080	)	,
(	13107	)	,
(	13133	)	,
(	13160	)	,
(	13186	)	,
(	13213	)	,
(	13240	)	,
(	13266	)	,
(	13293	)	,
(	13320	)	,
(	13347	)	,
(	13373	)	,
(	13400	)	,
(	13427	)	,
(	13454	)	,
(	13481	)	,
(	13508	)	,
(	13535	)	,
(	13562	)	,
(	13590	)	,
(	13617	)	,
(	13644	)	,
(	13671	)	,
(	13699	)	,
(	13726	)	,
(	13753	)	,
(	13781	)	,
(	13808	)	,
(	13836	)	,
(	13863	)	,
(	13891	)	,
(	13919	)	,
(	13946	)	,
(	13974	)	,
(	14002	)	,
(	14030	)	,
(	14058	)	,
(	14086	)	,
(	14114	)	,
(	14142	)	,
(	14170	)	,
(	14198	)	,
(	14226	)	,
(	14254	)	,
(	14282	)	,
(	14310	)	,
(	14339	)	,
(	14367	)	,
(	14395	)	,
(	14424	)	,
(	14452	)	,
(	14481	)	,
(	14509	)	,
(	14538	)	,
(	14567	)	,
(	14595	)	,
(	14624	)	,
(	14653	)	,
(	14681	)	,
(	14710	)	,
(	14739	)	,
(	14768	)	,
(	14797	)	,
(	14826	)	,
(	14855	)	,
(	14884	)	,
(	14913	)	,
(	14943	)	,
(	14972	)	,
(	15001	)	,
(	15030	)	,
(	15060	)	,
(	15089	)	,
(	15119	)	,
(	15148	)	,
(	15178	)	,
(	15207	)	,
(	15237	)	,
(	15266	)	,
(	15296	)	,
(	15326	)	,
(	15356	)	,
(	15386	)	,
(	15415	)	,
(	15445	)	,
(	15475	)	,
(	15505	)	,
(	15535	)	,
(	15566	)	,
(	15596	)	,
(	15626	)	,
(	15656	)	,
(	15686	)	,
(	15717	)	,
(	15747	)	,
(	15777	)	,
(	15808	)	,
(	15838	)	,
(	15869	)	,
(	15900	)	,
(	15930	)	,
(	15961	)	,
(	15992	)	,
(	16022	)	,
(	16053	)	,
(	16084	)	,
(	16115	)	,
(	16146	)	,
(	16177	)	,
(	16208	)	,
(	16239	)	,
(	16270	)	,
(	16301	)	,
(	16332	)	,
(	16364	)	,
(	16395	)	,
(	16426	)	,
(	16458	)	,
(	16489	)	,
(	16521	)	,
(	16552	)	,
(	16584	)	,
(	16615	)	,
(	16647	)	,
(	16679	)	,
(	16711	)	,
(	16742	)	,
(	16774	)	,
(	16806	)	,
(	16838	)	,
(	16870	)	,
(	16902	)	,
(	16934	)	,
(	16966	)	,
(	16998	)	,
(	17031	)	,
(	17063	)	,
(	17095	)	,
(	17128	)	,
(	17160	)	,
(	17192	)	,
(	17225	)	,
(	17257	)	,
(	17290	)	,
(	17323	)	,
(	17355	)	,
(	17388	)	,
(	17421	)	,
(	17454	)	,
(	17487	)	,
(	17519	)	,
(	17552	)	,
(	17585	)	,
(	17618	)	,
(	17652	)	,
(	17685	)	,
(	17718	)	,
(	17751	)	,
(	17784	)	,
(	17818	)	,
(	17851	)	,
(	17885	)	,
(	17918	)	,
(	17952	)	,
(	17985	)	,
(	18019	)	,
(	18052	)	,
(	18086	)	,
(	18120	)	,
(	18154	)	,
(	18188	)	,
(	18221	)	,
(	18255	)	,
(	18289	)	,
(	18323	)	,
(	18357	)	,
(	18392	)	,
(	18426	)	,
(	18460	)	,
(	18494	)	,
(	18529	)	,
(	18563	)	,
(	18597	)	,
(	18632	)	,
(	18666	)	,
(	18701	)	,
(	18736	)	,
(	18770	)	,
(	18805	)	,
(	18840	)	,
(	18875	)	,
(	18909	)	,
(	18944	)	,
(	18979	)	,
(	19014	)	,
(	19049	)	,
(	19084	)	,
(	19120	)	,
(	19155	)	,
(	19190	)	,
(	19225	)	,
(	19261	)	,
(	19296	)	,
(	19332	)	,
(	19367	)	,
(	19403	)	,
(	19438	)	,
(	19474	)	,
(	19510	)	,
(	19545	)	,
(	19581	)	,
(	19617	)	,
(	19653	)	,
(	19689	)	,
(	19725	)	,
(	19761	)	,
(	19797	)	,
(	19833	)	,
(	19869	)	,
(	19905	)	,
(	19942	)	,
(	19978	)	,
(	20014	)	,
(	20051	)	,
(	20087	)	,
(	20124	)	,
(	20160	)	,
(	20197	)	,
(	20234	)	,
(	20270	)	,
(	20307	)	,
(	20344	)	,
(	20381	)	,
(	20418	)	,
(	20455	)	,
(	20492	)	,
(	20529	)	,
(	20566	)	,
(	20603	)	,
(	20641	)	,
(	20678	)	,
(	20715	)	,
(	20753	)	,
(	20790	)	,
(	20828	)	,
(	20865	)	,
(	20903	)	,
(	20940	)	,
(	20978	)	,
(	21016	)	,
(	21054	)	,
(	21091	)	,
(	21129	)	,
(	21167	)	,
(	21205	)	,
(	21243	)	,
(	21281	)	,
(	21320	)	,
(	21358	)	,
(	21396	)	,
(	21434	)	,
(	21473	)	,
(	21511	)	,
(	21550	)	,
(	21588	)	,
(	21627	)	,
(	21665	)	,
(	21704	)	,
(	21743	)	,
(	21781	)	,
(	21820	)	,
(	21859	)	,
(	21898	)	,
(	21937	)	,
(	21976	)	,
(	22015	)	,
(	22054	)	,
(	22094	)	,
(	22133	)	,
(	22172	)	,
(	22211	)	,
(	22251	)	,
(	22290	)	,
(	22330	)	,
(	22369	)	,
(	22409	)	,
(	22449	)	,
(	22488	)	,
(	22528	)	,
(	22568	)	,
(	22608	)	,
(	22648	)	,
(	22688	)	,
(	22728	)	,
(	22768	)	,
(	22808	)	,
(	22848	)	,
(	22888	)	,
(	22929	)	,
(	22969	)	,
(	23010	)	,
(	23050	)	,
(	23091	)	,
(	23131	)	,
(	23172	)	,
(	23212	)	,
(	23253	)	,
(	23294	)	,
(	23335	)	,
(	23376	)	,
(	23417	)	,
(	23458	)	,
(	23499	)	,
(	23540	)	,
(	23581	)	,
(	23622	)	,
(	23663	)	,
(	23705	)	,
(	23746	)	,
(	23787	)	,
(	23829	)	,
(	23871	)	,
(	23912	)	,
(	23954	)	,
(	23995	)	,
(	24037	)	,
(	24079	)	,
(	24121	)	,
(	24163	)	,
(	24205	)	,
(	24247	)	,
(	24289	)	,
(	24331	)	,
(	24373	)	,
(	24416	)	,
(	24458	)	,
(	24500	)	,
(	24543	)	,
(	24585	)	,
(	24628	)	,
(	24670	)	,
(	24713	)	,
(	24756	)	,
(	24798	)	,
(	24841	)	,
(	24884	)	,
(	24927	)	,
(	24970	)	,
(	25013	)	,
(	25056	)	,
(	25099	)	,
(	25142	)	,
(	25185	)	,
(	25229	)	,
(	25272	)	,
(	25316	)	,
(	25359	)	,
(	25403	)	,
(	25446	)	,
(	25490	)	,
(	25533	)	,
(	25577	)	,
(	25621	)	,
(	25665	)	,
(	25709	)	,
(	25753	)	,
(	25797	)	,
(	25841	)	,
(	25885	)	,
(	25929	)	,
(	25974	)	,
(	26018	)	,
(	26062	)	,
(	26107	)	,
(	26151	)	,
(	26196	)	,
(	26240	)	,
(	26285	)	,
(	26330	)	,
(	26374	)	,
(	26419	)	,
(	26464	)	,
(	26509	)	,
(	26554	)	,
(	26599	)	,
(	26644	)	,
(	26689	)	,
(	26735	)	,
(	26780	)	,
(	26825	)	,
(	26871	)	,
(	26916	)	,
(	26962	)	,
(	27007	)	,
(	27053	)	,
(	27099	)	,
(	27144	)	,
(	27190	)	,
(	27236	)	,
(	27282	)	,
(	27328	)	,
(	27374	)	,
(	27420	)	,
(	27466	)	,
(	27513	)	,
(	27559	)	,
(	27605	)	,
(	27652	)	,
(	27698	)	,
(	27744	)	,
(	27791	)	,
(	27838	)	,
(	27884	)	,
(	27931	)	,
(	27978	)	,
(	28025	)	,
(	28072	)	,
(	28119	)	,
(	28166	)	,
(	28213	)	,
(	28260	)	,
(	28307	)	,
(	28354	)	,
(	28402	)	,
(	28449	)	,
(	28497	)	,
(	28544	)	,
(	28592	)	,
(	28639	)	,
(	28687	)	,
(	28735	)	,
(	28783	)	,
(	28830	)	,
(	28878	)	,
(	28926	)	,
(	28974	)	,
(	29023	)	,
(	29071	)	,
(	29119	)	,
(	29167	)	,
(	29216	)	,
(	29264	)	,
(	29312	)	,
(	29361	)	,
(	29410	)	,
(	29458	)	,
(	29507	)	,
(	29556	)	,
(	29604	)	,
(	29653	)	,
(	29702	)	,
(	29751	)	,
(	29800	)	,
(	29850	)	,
(	29899	)	,
(	29948	)	,
(	29997	)	,
(	30047	)	,
(	30096	)	,
(	30146	)	,
(	30195	)	,
(	30245	)	,
(	30294	)	,
(	30344	)	,
(	30394	)	,
(	30444	)	,
(	30494	)	,
(	30544	)	,
(	30594	)	,
(	30644	)	,
(	30694	)	,
(	30744	)	,
(	30795	)	,
(	30845	)	,
(	30895	)	,
(	30946	)	,
(	30996	)	,
(	31047	)	,
(	31098	)	,
(	31148	)	,
(	31199	)	,
(	31250	)	,
(	31301	)	,
(	31352	)	,
(	31403	)	,
(	31454	)	,
(	31505	)	,
(	31557	)	,
(	31608	)	,
(	31659	)	,
(	31711	)	,
(	31762	)	,
(	31814	)	,
(	31865	)	,
(	31917	)	,
(	31969	)	,
(	32020	)	,
(	32072	)	,
(	32124	)	,
(	32176	)	,
(	32228	)	,
(	32280	)	,
(	32332	)	,
(	32385	)	,
(	32437	)	,
(	32489	)	,
(	32542	)	,
(	32594	)	,
(	32647	)	,
(	32699	)	,
(	32752	)	,
(	32805	)	,
(	32858	)	,
(	32911	)	,
(	32963	)	,
(	33016	)	,
(	33070	)	,
(	33123	)	,
(	33176	)	,
(	33229	)	,
(	33282	)	,
(	33336	)	,
(	33389	)	,
(	33443	)	,
(	33496	)	,
(	33550	)	,
(	33604	)	,
(	33657	)	,
(	33711	)	,
(	33765	)	,
(	33819	)	,
(	33873	)	,
(	33927	)	,
(	33981	)	,
(	34036	)	,
(	34090	)	,
(	34144	)	,
(	34199	)	,
(	34253	)	,
(	34308	)	,
(	34362	)	,
(	34417	)	,
(	34472	)	,
(	34526	)	,
(	34581	)	,
(	34636	)	,
(	34691	)	,
(	34746	)	,
(	34801	)	,
(	34857	)	,
(	34912	)	,
(	34967	)	,
(	35023	)	,
(	35078	)	,
(	35134	)	,
(	35189	)	,
(	35245	)	,
(	35301	)	,
(	35356	)	,
(	35412	)	,
(	35468	)	,
(	35524	)	,
(	35580	)	,
(	35636	)	,
(	35692	)	,
(	35749	)	,
(	35805	)	,
(	35861	)	,
(	35918	)	,
(	35974	)	,
(	36031	)	,
(	36088	)	,
(	36144	)	,
(	36201	)	,
(	36258	)	,
(	36315	)	,
(	36372	)	,
(	36429	)	,
(	36486	)	,
(	36543	)	,
(	36600	)	,
(	36658	)	,
(	36715	)	,
(	36773	)	,
(	36830	)	,
(	36888	)	,
(	36945	)	,
(	37003	)	,
(	37061	)	,
(	37119	)	,
(	37177	)	,
(	37235	)	,
(	37293	)	,
(	37351	)	,
(	37409	)	,
(	37467	)	,
(	37526	)	,
(	37584	)	,
(	37643	)	,
(	37701	)	,
(	37760	)	,
(	37818	)	,
(	37877	)	,
(	37936	)	,
(	37995	)	,
(	38054	)	,
(	38113	)	,
(	38172	)	,
(	38231	)	,
(	38290	)	,
(	38350	)	,
(	38409	)	,
(	38468	)	,
(	38528	)	,
(	38587	)	,
(	38647	)	,
(	38707	)	,
(	38767	)	,
(	38826	)	,
(	38886	)	,
(	38946	)	,
(	39006	)	,
(	39066	)	,
(	39127	)	,
(	39187	)	,
(	39247	)	,
(	39308	)	,
(	39368	)	,
(	39429	)	,
(	39489	)	,
(	39550	)	,
(	39611	)	,
(	39671	)	,
(	39732	)	,
(	39793	)	,
(	39854	)	,
(	39915	)	,
(	39977	)	,
(	40038	)	,
(	40099	)	,
(	40161	)	,
(	40222	)	,
(	40283	)	,
(	40345	)	,
(	40407	)	,
(	40468	)	,
(	40530	)	,
(	40592	)	,
(	40654	)	,
(	40716	)	,
(	40778	)	,
(	40840	)	,
(	40903	)	,
(	40965	)	,
(	41027	)	,
(	41090	)	,
(	41152	)	,
(	41215	)	,
(	41277	)	,
(	41340	)	,
(	41403	)	,
(	41466	)	,
(	41529	)	,
(	41592	)	,
(	41655	)	,
(	41718	)	,
(	41781	)	,
(	41845	)		 -- array index 4095 (voltage = "111111111111" or 4095 mV), distance output 3787 (37.87 cm)

);


end package LUT_pkg;
